// ram_write.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ram_write_tb (
		//input  wire        clk_clk,                                //             clk.clk
		//input  wire [31:0] ram_w_0_control_control_write_base,     // ram_w_0_control.control_write_base
		//input  wire [31:0] ram_w_0_control_control_write_length,   //                .control_write_length
		//output wire        ram_w_0_control_control_done,           //                .control_done
		//input  wire        ram_w_0_control_control_fixed_location, //                .control_fixed_location
		//input  wire        ram_w_0_control_control_go,             //                .control_go
		//input  wire        ram_w_0_user_user_write_buffer,         //    ram_w_0_user.user_write_buffer
		//input  wire [31:0] ram_w_0_user_user_buffer_data,          //                .user_buffer_data
		//output wire        ram_w_0_user_user_buffer_full,          //                .user_buffer_full
		//input  wire        reset_reset_n                           //           reset.reset_n
	);

	reg          clk_clk = 1'b0;
        reg          reset_reset_n = 1'b1;
        // Declare input signals as reg
        reg [31:0] ram_w_0_control_control_write_base;
        reg [31:0] ram_w_0_control_control_write_length;
        reg        ram_w_0_control_control_go;
	wire       ram_w_0_control_control_done;
	reg        ram_w_0_control_control_fixed_location;
        reg [31:0] ram_w_0_user_user_buffer_data;
        reg        ram_w_0_user_user_write_buffer;
	wire       ram_w_0_user_user_buffer_full;

	wire         ram_w_0_avalon_master_waitrequest;                // mm_interconnect_0:ram_w_0_avalon_master_waitrequest -> ram_w_0:M_AVALON_WAITREQUEST
	wire  [31:0] ram_w_0_avalon_master_address;                    // ram_w_0:M_AVALON_ADDRESS -> mm_interconnect_0:ram_w_0_avalon_master_address
	wire   [3:0] ram_w_0_avalon_master_byteenable;                 // ram_w_0:M_AVALON_BYTEENABLE -> mm_interconnect_0:ram_w_0_avalon_master_byteenable
	wire         ram_w_0_avalon_master_write;                      // ram_w_0:M_AVALON_WRITE -> mm_interconnect_0:ram_w_0_avalon_master_write
	wire  [31:0] ram_w_0_avalon_master_writedata;                  // ram_w_0:M_AVALON_WRITEDATA -> mm_interconnect_0:ram_w_0_avalon_master_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect; // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s1_address;    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable; // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [mm_interconnect_0:ram_w_0_reset_sink_reset_bridge_in_reset_reset, onchip_memory2_0:reset, ram_w_0:M_AVALON_RSTN]

	localparam  CLOCK_PERIOD            = 10; // Clock period in ps
        localparam  INITIAL_RESET_CYCLES    = 1000;  // Number of cycles to reset when simulation starts

	ram_write_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (1'b0),                                             // (terminated)
		.freeze     (1'b0)                                              // (terminated)
	);

	write_ram #(
		.AVALON_DATA_WIDTH    (32),
		.FIFO_DEPTH           (4),
		.FIFO_DEPTH_LOG2      (2),
		.AVALON_ADDRESS_WIDTH (32)
	) ram_w_0 (
		.control_write_base     (ram_w_0_control_control_write_base),     //       control.control_write_base
		.control_write_length   (ram_w_0_control_control_write_length),   //              .control_write_length
		.control_done           (ram_w_0_control_control_done),           //              .control_done
		.control_fixed_location (ram_w_0_control_control_fixed_location), //              .control_fixed_location
		.control_go             (ram_w_0_control_control_go),             //              .control_go
		.user_write_buffer      (ram_w_0_user_user_write_buffer),         //          user.user_write_buffer
		.user_buffer_data       (ram_w_0_user_user_buffer_data),          //              .user_buffer_data
		.user_buffer_full       (ram_w_0_user_user_buffer_full),          //              .user_buffer_full
		.M_AVALON_WAITREQUEST   (ram_w_0_avalon_master_waitrequest),      // avalon_master.waitrequest
		.M_AVALON_ADDRESS       (ram_w_0_avalon_master_address),          //              .address
		.M_AVALON_WRITE         (ram_w_0_avalon_master_write),            //              .write
		.M_AVALON_BYTEENABLE    (ram_w_0_avalon_master_byteenable),       //              .byteenable
		.M_AVALON_WRITEDATA     (ram_w_0_avalon_master_writedata),        //              .writedata
		.M_AVALON_CLK           (clk_clk),                                //    clock_sink.clk
		.M_AVALON_RSTN          (~rst_controller_reset_out_reset)         //    reset_sink.reset_n
	);

	ram_write_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                          //                                clk_0_clk.clk
		.ram_w_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // ram_w_0_reset_sink_reset_bridge_in_reset.reset
		.ram_w_0_avalon_master_address                  (ram_w_0_avalon_master_address),                    //                    ram_w_0_avalon_master.address
		.ram_w_0_avalon_master_waitrequest              (ram_w_0_avalon_master_waitrequest),                //                                         .waitrequest
		.ram_w_0_avalon_master_byteenable               (ram_w_0_avalon_master_byteenable),                 //                                         .byteenable
		.ram_w_0_avalon_master_write                    (ram_w_0_avalon_master_write),                      //                                         .write
		.ram_w_0_avalon_master_writedata                (ram_w_0_avalon_master_writedata),                  //                                         .writedata
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),    //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                         .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	// Clock signal generator
   always begin
      #(CLOCK_PERIOD / 2);
      clk_clk = ~clk_clk;
   end
   
   // Initial reset
   initial begin
      //repeat(INITIAL_RESET_CYCLES) @(posedge clk_clk);
      #0 
      reset_reset_n = 1'b0;
      #20; reset_reset_n = 1'b1; 
   end
	integer i;
	parameter TOGGLE_CYCLES = 10;
  // Stimulus for the testbench
    initial begin
        // Wait for the reset de-assertion

        // Initialize inputs
        ram_w_0_control_control_write_base = 32'h00000000;
        ram_w_0_control_control_write_length = 32'h0000000C;
        ram_w_0_control_control_go = 1'b0;
	ram_w_0_control_control_fixed_location = 1'b0;
        ram_w_0_user_user_buffer_data = 32'hA5A5A5A5;
        ram_w_0_user_user_write_buffer = 1'b0;

        // Wait for a few clock cycles
        repeat(2) @(posedge clk_clk);
	end

        // Trigger the input signals
	initial begin
        #0
        ram_w_0_user_user_write_buffer = 1'b1;
        wait (ram_w_0_user_user_buffer_full)
	ram_w_0_user_user_write_buffer = 1'b0;
        end

	initial begin
	#195
    // Infinite loop
    forever begin
        // Set control signal to 1
	wait (ram_w_0_control_control_done);
        ram_w_0_control_control_go = 1;
        
        // Wait for 5 time units
        #5;
        
        // Set control signal to 0
        ram_w_0_control_control_go = 0;
        
        // Wait for 5 time units
        //#20;
    end
end
    
	initial begin
	// Trigger the input signals
        #400
	ram_w_0_control_control_fixed_location = 1'b1;
        #600
        $finish;
    end

endmodule
